/*
*
* Copyright 2023 Massimo Vincenzi
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*    http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
*/
`ifndef SV_APB_SEQUENCER
`define SV_APB_SEQUENCER

class apb_sequencer extends uvm_sequencer #(apb_trans_item, apb_trans_item);
	`uvm_component_utils(apb_sequencer)

	function new(string name = "apb_sequencer", uvm_component parent = null);
		super.new(name, parent);
	endfunction

endclass : apb_sequencer

`endif